class apb_gen;
	// Constructor
	function new();
	endfunction

	// Run task
	task run();
		$display("### Inside run task of generator");
	endtask
endclass
