class apb_bfm;
	// Constructor
	function new();
	endfunction

	// Run task
	task run();
		$display("### Inside run task of bfm");
	endtask
endclass
