`include "apb_common.sv"
`include "apb.v"
`include "mem.v"
`include "apb_intf.sv"
`include "apb_tx.sv"
`include "apb_gen.sv"
`include "apb_bfm.sv"
`include "apb_mon.sv"
`include "apb_cov.sv"
`include "apb_agent.sv"
`include "apb_sbd.sv"
`include "apb_env.sv"
`include "top.sv"
