class apb_cov;
	// Constructor
	function new();
	endfunction

	// Run task
	task run();
		$display("### Inside run task of coverage");
	endtask
endclass
