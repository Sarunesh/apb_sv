class apb_sbd;
	// Constructor
	function new();
	endfunction

	// Run task
	task run();
		$display("### Inside run task of scoreboard");
	endtask
endclass
