class apb_mon;
	// Constructor
	function new();
	endfunction

	// Run task
	task run();
		$display("### Inside run task of monitor");
	endtask
endclass
